module moduleName #(
parameter
) (
input wire              i_ref_clk;
input wire              i_rst_n;
input wire              i_clk_en;
input wire              i_div_ratio;
output reg              o_div_clk;            
);
    
endmodule